// `timescale  1ns / 1ns

//----------------------------------------------------------------
// Declare
//----------------------------------------------------------------

// This Template is written by Pu Junhao, which you can adjusted depending on your own style.
// Declare your information here.
// You may wanna use UTF-8. Delcare it here.
// You may wanna declare copyrights here. ALL RIGHTS RESERVED BY PU JUNHAO.

module code

//----------------------------------------------------------------
// Inherited Module Params
//----------------------------------------------------------------

#(
    parameter PARAM = 0
)

//----------------------------------------------------------------
// Ports
//----------------------------------------------------------------

(
     clk_i
    ,rst_i
    ,out_o
);

    // Inputs
    input clk_i;
    input rst_i;

    // Outputs
    output reg [31:0] out_o;

//----------------------------------------------------------------
// Registers / Wires / Params / Includes
//----------------------------------------------------------------

// `include "defs.v"
localparam
    PARAM1 = 1,
    PARAM2 = 2;

reg [31:0] ROM[255:0]; //31x256
reg [31:0] state;
reg [31:0] state_cnt;

wire state_pulse;

integer row;

genvar gen_row;

//----------------------------------------------------------------
// Test Bench
//----------------------------------------------------------------

// // Uncommenting This Part First

// // code Parameters
// parameter PERIOD = 10;

// // code Inputs
// reg   clk_i = 0;
// reg   rst_i = 0;

// // code Outputs
// wire  [31:0]  out_o;    

// initial begin
//     forever #(PERIOD/2)  clk_i = ~ clk_i;
// end

// initial begin
//     #(PERIOD*2) rst_i  =  1;
// end

// initial begin
//     // Write Test Bench Here
//     $finish;
// end

//----------------------------------------------------------------
// Circuits
//----------------------------------------------------------------

// Initialization
initial begin
    for(row = 0; row <= 255; row = row + 1)
        row = row + 1;
end

// State Machine
always @(posedge clk_i) begin
    if (rst_i == 1) begin
        row = 0;
    end
    else begin
        row = row + 1;
    end
end

endmodule


//----------------------------------------------------------------
// Personalized label
//----------------------------------------------------------------

// Keep your own style!

// OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOoooo**.........*..*.  ......*********,ooooooooooooooooooooooooooOOOOOOOO\*[oooO@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@OooOO@OO@@@OO@@@OOOOOOOOO@@OO^...
// OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOooooo`*******..........     .....*********\oooooooooooooooooooo[`***,\OOOOOOOO\*.,O@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@OO@@@O@@@@@@@@@@@@@@@OOOOOO^...
// OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOoo`***.................   .....*****************************************,\OOO@@@OO\*O@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@OOO@O@@@@@@o\O@@@@@@@O^...
// OOOOOOOOOOOOOOOOOOOOOOOOOOOOOoooo]**...................   .*,]]***********************,]]oOOOOOOOOOOo]]]*=OOOOOOOOOO/O@@@@@@@@@@@@@@@@@@@@@@@@@OOO@@@@@@@@@@@@OOOO\O@@@@@@@@@@O^...
// *****************=oOOOOOOOOOOOOOooo^*******]]]*******....**]O@@@OOO\`************,/oOOOOOOOOOOOOOOOOOOOOOOOOOOoOOOOo]o@@@@@@@@@@@@@@@@@OOOOOOOOOOO@@@@@@@@@@@@@OO@OOOOOOOOOOO@O^***
// OOOOOOOOOOOOOOOOo=OOOOOOOOOOOOOOooo***************[****=*.=OOOOO@@@@@OOo]**]ooOOOOOoOOOOOOOOOOooooooo/[[[\oOOOOOO@@@@@@@@@@@@@@@@@OO@@@OOOOOOOOOOO@@@@@OOOO@@@@@@@@@@@@@@@@@@@O^**`
// OOOOO@@@@OOO@@@Oo=OOOOOOOOOOOOOooooo/*..............**o`..........[OO@@@@OOo[\OOOoooooOOOOOOOOOO\*............=O@@@@@@@@@@@@@@@@@OOoO@@@OOOoooOOOO@@@OOOOOOOOO@@@@@@@@@@@@@@@@Ooooo
// OOOOO@@@@OOO@@@Oo=OOOOOOOOOOoooo[`**...................       ..*]]/oO@@@@@@^*[[...            ...,\OO\`......,O@@@@@@@@@@@@@@@@@OOOoO@@@@Oo*=ooooOOOooooOOO/[\O@@@@@@@@@@@@@@OOooo
// O@@OO@@@@@OO@@@OO=OOOOOOOOoo`****..................             .,@@OO@@@@@@O^.                       .,OOOooooooO@@@@@@@@@@@@@@@@OOo,@@@@@^**[/[/\oooooo/*.....=O@@@@@@@@@@@@OOOoo
// O@@OO@@@@@OO@@@@O*oOOOOOoo`*..........**,ooo/`.              ../OOoooOOO[[..........                      .,\OOOoOOO@@@@@@@@@@@@@@@OOOO@@@@O*.*****o/*,/o`....*=OO@@@@@@@@@@OOOOooo
// O@@OOO@@@OOOOOOOO*oOOOOo/*..........**/oOOO`.       .   .  ./Ooooo`.//....................                    .[OOOOOO@@@@@@@@@@@@@@@@@@@@@@O`..,OO`*=oO@O...*/OOO@@@@@@@@@OOOOoooo
// O@@OOOOOOOoOOOOOOooOOOOo^*.......*/oooOOO`         ..   .,Oo[,o/...,...............*..........                   ,\O@@@@@@@@@@@@@@@@@@O/`\O@@@@@@@@/*.*,[`**,oOOOOO@@@@@@@@Oooooooo
// O@@OO@@@@@OO@@`.,[OOOOOoo*......*=ooOOOOo.         ..   ,[`*,o.. ..............    ..............           ..     .[oO@@@@@@@OO@@@@@@O\]/O@@@@@@@@O\]*.***,oOOOOOOO@@@@@@@@OOooooo
// O@@OOO@@@OOO@^.......[OOOO\.....*=oOO@OOo.        ...   .****.  ................       ...      ....         ..     ...,O@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@O`*/ooOOOOOOO@@@@@@OOOOooooo
// OO@OOOOOOOOOO............,[Oo]*.*=O@@OOOO^.     .,O@^....=`.... ...............*..                 ...                ....\@@@@@@@@@@@@@@O@@@@@@\/@@@@@@O]OOOOOOOOOO@@@@@@OooOOo***
// OO@OO@@@@@O@^................,OOO@@@OOOOOO`..,]/O@OOO`............   ....... ..*....                  ..             .......O@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@OOo\/OOo`*
// O@@OOO@O@OOO`...........*....*/O@@@@@@OOOOOOOO@@OOOO`=`....=O^...         ..  .......                                    ....,O@@@@@@@@@@O@@@@@@@@@@@OOOO@@@@@@@@@@@@@@@@@OOOOOOOOO
// O@@OOOOOOOO/..........*]]]]]O@@@@@@@@@@@OOOO@@@OOOO^..=\...**. ..         ..  .  ..               .                        ....,@@@@@@@@@O@@@@@@@@@@O`**oOOO@@@@@@@@@@@@OOooOO^....
// OO@OO@@@@@O^........,ooOOOOO@@@@@OO[\O@@@@@@@OOOO/`....,o\`***..          .   .   ..   .....        ..                      ..  .\@@@@@@@@@@@@@@@@@@O\***oOOOOOO@@@OooOOOo\**......
// OO@OOO@O@@O.......*/Oo*.*O@@@@@Oo*..*=@@@@@OOOO/.........=OO\`**..        .  ..   ...          .    ...........               .. .,O@@@@@@@@@@@@@@@@@@O\]oOOOOOOO@@@@OOooo/*.*****.
// O@@OOOOOO@^......*oOO^...=@@@@@OOO\]/@@@@@OOO`...........=@@@Oo]/\..      .  ..    ..          ..........*]**..                ..  .\@@@@@@@@@@@@@@@@@@OOOOOOOO@@@@@@@@@Ooooooooooo
// O@@OO@@@@O^.....,oOOOooooOO@@@@OOO@@@@@@OOO^........... .O@@O....****... ..   .    ...          ........*o^*,`*..         ....  ... .,O@@@@@@@@@@@@@@@@@O@@@@@@@@@@@@@@@@@O\]]/oooo
// OO@OOO@@@O*.....=oOOOOOOO/*,O@@@OOO@@@@OOO`..... .....  =@O[*.   ..............     ..            ......*.,oOO^*.         ..o`.,OO.   .\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@OO
// O@@OOOOO@^......*\OOOOOOOO...\@OO@@@@OOO/. .. ..  ..   .OO`...    ..     ..   .      .             .......*[[[`*.        ..*[`..=Oo.   .=@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@O\..
// O@@OO@@@@^.......*[[*[OOOO`*.,OO]O@@OOO^.  .. .. ..    =O^....     ..    ..   .                     ...**.,OO^*............*..=oOoo].    ,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@O^..[OO
// OO@OOOO@O^...**.**.....=OOOOooO@@@@OOO`.   .. .....   .=/.  ..     ...   ..   .                         ......*....**.....**..,o^*\OOO`. .=@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@`...[\OO\]
// OO@OOOOOO^....******.*/oooOOOOO@@OOOO`.   ..  ....    .=`   ...     ..   ..   .                            ..*^*........**.*=o[**/OO@@@O. .=@@@@@@@@@@@@@@@@@@@@@@@@@@@O[oo]....,\O
// OO@OO@@@O^....******=ooOO/[[\O@@OOOO^.    ... ....    ...    ..      ... ..    .    .                        .*........**...   ,oOO@@@@@O. .OOO@@@@@@@@@@@@@@@@@@@@@@@@OOO`*[\O\].,
// OO@OOOO@OOOOOOOooooOO@@@@OOOO@@OOOOO.     ........     .      ...     .....         ..      ..         .      .......,o\*...../OOO@@@@@@@\. .OO@@@@@@@O@@@@@@@@@@@@@@@O`*\O@O`..,\@
// OO@OOOOOOOOOOO@@@@@@@@@@@@@@@@OOOOO`      ........             ...    .....         ..       .  .              .,OOOoooooooOOOOOO@@OO@@@@@^ .=@OOO`.O^.O@@@@@@@@OOO@@O..[O\`,\O\]/O
// OO@OO@@@@@OOOO@OOO@@@@@@@@@@OOOOO@/.      ........     ....      ...  .....         ..       .. ..       .      .=ooooOOOOOOO@@@@@@@@@@@@O`  .O\O^.=O*.o`,@@@@@@@OOOOOOO`..[OO`,O@O
// O@@O/....OOOO@O^..*OOO@@@@@OOO`*OO..      .........    ......     =O`........       ...      ..  ....    ...    ..=ooOO@OOOOO@@@/\O@@@@OO.    *OO..OO*=O..O/.\@@@OOOOOOOOOO`.,OO@@@
// @OOOO....OOO@@OO`*/OOOO@@@OO`..OO`.       ..........    .    .    .O/o`.......      ...      .\.  ...........    ..=oO@@@@@@@@O`*.*]oOOOO^.   .O\.,O^*OO.=O^.=OOO/oOOOOOOOOOOOoO@OO
// O@OOOOOOOOO@@@@@@@@@@@@@@O/.,/@@^.....    ...........         ... .,*..**.......     ..      .*... ............   ..\O@@@@@@[...*/OOOOOOO^.    =O,Oo.=O^./O../OOo/oOOOOOOOOOOoOO@@O
// O@@OOOOOOOOO@@@@@@@@@@@@/,]oO@@^......     ...........             ...  ...**...*..  ..      .*.... .................\OOO/`..*.*oOOOo*\OO^.    .OOO^.=O..OO..OOOO^=O@@OOOO[*.,ooOOO
// O@@@@OOOO@@@@@@@@@@@@@@OooOO@@O........   ...*.........             ..   .. ..******..*. ..  .*........o`.............,[.  .=^./OO/*\oOOO^     .\@@^.o/.=O^..OOOO^*O@@@OOOOOOooOooO
// O@@OO@@@@@@@@@@@@@@@@@/[[O@@@@O..... ... .............*.             ..  ..     ....*\O\]].  ..... ......**............**. .=..OOOO\oOOOO^     .,@@OOO^./@^.=@@OOo*oOOOOOOO^**,o`..
// O@@OO@@@@@@@@@@@@@@@O.  .O@@O@/.....   ..  ..............             .  ..          .,*,[.  .....    ..*....**o\]]*....*.  =*.OOOOO*.OOO.     ..O@@@@\/@@`,/@@@OooOO@@@OOO^=o\,o`.
// O@@OOO@@@@@@@@@@@@@@`  ,@@@OO@` ...     .  ...............            ......         .*....  ..............**..**[OO\*..**. .=*,OOOOOOOOO.     ..OOOOO@@@@@@@@@@OOOOO@OOOo`**[[*=^.
// O@@OO@@@@@@@@@@@@@@^. ,O@@@O@O. ...     .. .................           ......        .*....   .........     ...****,[\^*.*.. .,**oOOOOOOO.     ..O@OO@@@@@@@@OOOoOOOOOOOO\*.*,]`=^.
// O@@OO@@@@@@@@@@@@@@. ,O@@@OO@`  ...        ... ...*.    .......         ...*.        .*....  ....*/*.. ... .............=\`.   ..*\oooOOO.    ...O@O@@@@@@@OOOOOOOOOOO@OOOOO]*..,`.
// O@@OOO@@@OOO@@@@@@/.,O@@@@O@O.   ..        ...  ..\^.    .=*.........   ....o.       .*........***..............      ...=O\.     ....,O..    . .=@@@@@@@@@OOOOOOOOOOOOOOOOOOo]`...
// O@@OO@@@@@O@@@@@@@`.O@@@@@O@^    ..        .*.   .=o.     .,`........    ..*O\.      .*....***=[...............        ...,O\.         ........  =@O@@@@@@@OOOOOOOOOOOOOoo\/OOO^...
// O@@OO@@@@@O@@@O@@O./@@@@@OOO.    ..        .o^   .=/\.     .,\*.............=@^.    ..*../OOOo***..........       .......,.=O^   .     ........  .OoO@@@@@@@@O@@OOOOOOOOOOooo[`*...
// O@@OO@@@@@@@@@@@@^=@@@@@@oO^      .        .\\.  .=^....  ....****..........,OO`.   ...,OOo*....................]]OO@@@@/...\O`  ..    .......   .OO/o@@@@@OOO@@OooOOOo[**.......]O
// O@@OO@@@@@@@@@@@@\@@@@@@@OO. .     .       .O@.   .*..............***........,OO`.  ..*[.=o..........*,]]/OOOOO@@@@@@@O`.....O^ ...    .*....    .OO^*\@@@@@OOOO`oO\*\^.......,OOOO
// O@@OO@@@@@@@@@@@.=@@@@@@@O....     .     ...O@^   .*............*]...*[o]`....=OO....*...=o....*]]OOO@OOOO/......\O/\@/......=\....   .,*...     .O@O^=O@@OO^....,`*..`*..........*
// O@@@@@@@@@@@@@O..@@@@@@@@@`...     ..  ....,O@O.....*............,O^.....*[\`*]]/[[\o^**,oo../@@@@@O^............=O^.........,O..... ..o`..      .=OOooO@O]......,oo..**...........
// O@@@@@@@@@@@@O..O@@@@@@@@@^.,*      .......=OOO^....*.....  .......\O`.........*OOOoooo\]]*..[[....o^............=O^..........O........O.         =OOooO@@@OO]oooOo*.,\*]]]]]]O\OOO
// @@@@@@@@@@@@O. =@@@@@@@@@@^..*.     .......=OO`.....................,\o`*.......*oOO***oO/....    .,/......     .=^...........=*.*.........    .. =OOOoO@@@@@OOOOOOOOOOOO@@@@@@@OO.
// @@@@@@@@@@@@^. =O@OOOO@@@@^ ....    .......=OO..,]***ooooooOOO/`.......**``*...***[***=OO.....     ......     ..=`............=^.**.......     .. =@@@OO@@@OOOOOOOOOOOOOOOOO@OOOOO\
// O@@@@@@@@@@@^. =O@@OOOO@@@^..O*...   ......=O^.......*,[[`/*....     ....******.*****,OOo......     ..,o]...,]o`..............=^*....=O^.      .*.=@@@OO@@OOOOOOOOOOOOOOOOOOOOooooO
// O@@OO@@@@@@@^. =OOO@OoO@@@^..O^...*........=O^.......................       .,OO\****\O`*[*.....     .........................=*..**,oO.      ..O.=O/\OOOOoO,OOOOooooooOOOOOOOOOOOO
// O@@OO@@@@@O@@`..OOO@@OO@@@\..OO.      .*...=O^...............,oOOOO\..       ...**]]**\OO`........    ........................Oo***,ooo...    .=@^=o,O@OOO=^.=OOOOOOOooooOOOOO@OO@O
// O@@OO@@@@OOO@O`.OO@@@@@@@@O..=@^.      .*..=OO..........,OOOOOO/[[[[^.   ....***...,OO`.,oOo]]]`**...........................=O/**/O/o...     .=O^=OO@OOOO*^..o[^,\OOooooooOOOO@@@@
// O@@OO@@@@@O@@OOO`=@OO@@@@@@^.=@@`.     ..***O@^.....,/@@@OO[........*..  ......   ....**.....................................O/***[`**...     .OO^=O@OOOOo*^..***...,\oooooOOOoO@@@
// O@@OO@@@@OO@OOO@OOOOO@@@@@@O..O@@\.     .***O@O..,/@@@OO@\...........*.         ....  ..**.......  ........................./O^.....,...      .OO*=O@OOOO^*^..*........[[ooOOo*.\O@
// O@@OO@@@@@@@OOO@O@@O@@@@@@@@O.=@@@\..    .**\@@O,\@@@@O.,O\......   ....                ..*`.  ............................=O^.....,`...     .=OO*=O@@@@O**^..*............*\o...=O
// O@@OO@@@@@@OOO@@@@@@@@@@@@@O@\*O@@@\..    .^=@@@O....,O\.......    .*...                   ....    .......................,O`./o...,....     .O@O^=O@@@@O.=^..**....  ..   ........
// O@@OO@@@@@@OOO@@@@@@@@@@@@`=@@\*O@@@\..    ,oO@@@O..........,\o]]]//....                          .......................*..,OO^........    ..O@O^*O@@@@O.o^..*^.....        .... .
// O@@OO@@@@@@@@@@@@@@@@@@@@`.=@@@@OO@@@\..    .O@@@@@`......................   ..                    ..........................o/........   ...=O@O`*O@@@@^*o^..*^.  ..         .....
// O@@OO@@@@@@@@@@@@@@@@@@@^..=@@@OOOOO@@O`.    .O@OOOO....................... ...                     ........................*[.........  ....=O@o**O@@@O*.*^..*^.  ...         ....
// O@@OO@@@@@@@@@@@@@@@@@@/....@@O`,O@@@@@^......,O@OOO^..........................                      .......................,.........  ....*O@@^*=O@@@o`..^..*^.   ...        ....
// O@@OO@@@@@@@@@@@@@@@@@@^....O@O**,O@@@/[oO\`...,O@@@O^......................                         ......   .............,o**.............=O@@^*oO@@Oo^..*..*^.    ...        .=`
// O@@OO@@@@@@@@@@@@@@@@@@... .=@O*..=OOOO...,OO`...,OO@@\......................                         .....................Oo*..............oO@O^,O@OOoO^.....*^.     ..        .=o
// O@@O@@@@@@@@@@@@@@@@@@@^.  .=Oo*..=O@/\\...,\Oo*...\@@@\......................                            ................/O`..............=OO@O`=@OOo=O*.....*^.      ..       ..\
// O@@@@@@@@@@@@@@@@@@@@@@O.  ..O/*..=O@O**^......=OO`..[@@O.....................                           .       ........//................OO@@^=@OOO`OO......=^.       ..       ..
// O@@@@@@@@@@@@@@@@@@@@@@@\. ..o^...*O@*o`.......=@@@@@O`.,o\..................                                     ......*..........*....../OO@O*OOOO^*O^......=^.        ..      ..
// O@@@@@@@@@@@@@@@@@@@@@@@@^. .\o*..=O@..*`.......\@@@@@@@@@O/`**..............         .....       ..            .................**......=@@OO*=OOOO*=O`......o\.        ...     ..
// @O@@@@@@@@@@@@@@@@@@@@@@@O`..=O*.=O@@^..**........\@@@@@@@@\.................        .......                    ............,]O^**......,@@O/*/OOOO^./O......,Oo.    ..   ...     .
// O@@O@@@@@@@@@@@@@@@@@OO/..=...O`.\@@@O. ..\.........\@@@@@@@\...............          ..                     ....***.....]/O@@O`*...o...OO`*/OOOOOO`*OO.... .=O^..    .    ...    .
// @@O@@@@@@@@@@@@@@@@/......=O..\O^*O@OO^.  .O\....*....,O@@@@@O`..........                                  ...**..*....=oooo@@^....=o...*]O@@OOOOOo*/O^......=O*..    ..    ...    
// OOO@@@@@@@@@@@@@@@/.  ....O@\.,OOO@@OOO`. ..O@\.  ..O@@@OO@@@@@^........                                      ........*****o@/....=@Oo@@@@@@@OOOOO/*OO^......oo*..     ..    ...   
// OO@@@@@OO/`*O@@@@O.. .....OOO^.O@@@O.OOO....=@@@\.   .,@@@O`[O@@O`...                                       .......********oO`....O@OO@@@@@@@@OOOO^=OO*....../**...    ..     ...  
// O@@@Oo`.. .=O@@@O`.......=O@@@\*O@@^.,OOO...=@@@@@O`.  .,O@O^.,O@@@\..                                  .........***********...../OO@@@@@@@@@@OOOO*oOO*.......**...     ..     ....
// @@O/..    ,O@@@^.........OO@@@@O`\O...=OO\..=@@@@@@@@O`. ..[`.  .\@@@@\`..                        .............************...../OO@@@@@@@@@@@OOOO*OOO^........*...     ...     ...
// @O/..   .,O@@@@..........OO@@@@@OO\*. .=OO^.=@@@@@@@@@@@O\].,..   ,O@O@@@OO]...               .............***************...../@O@@@@@@@@@@@@@OO/*OOO^....]........     ..     ...
// O\*..  .,@@@@@/.........=OO@O@@@@@O.*]..OO`.=@@@@@@@@@@@@@@@@O^.   ,OOOOOOOOOOOOO]]]....................,]o`*]************...*O@OOO@@@@@@@@@@@@OOo,OOO^.../O^.......     ...     ..
// o/..  .,O@@@@@^.........OOO@@@@@@@^  ..*,`..=@@@@@@@@@@@@@@@@@@^.   .\OOOOOOOOOOOO@@@@OOO\]]]]]]..*]]ooooooooooooo]***,oo`*.,OOOOOO@@@@@@@@@@@@@OO*OOO.../OOo.......      ...     .
// o... .,O@@@@@@^........=OOO@@@@@@O.     ....=@@@@@@@@@@@@@@@@O/o.    .**...,[OO@@OOOOoOO@@@@@@@@@OOOOooooooooooooooo*ooo`..*ooOOOOO@@@@@@@@@@@@@OO*OOO...OOOO^.......     ...      
// *....=O@OO@@@O.........oO/o@@@@@@^.    .....=@@@@@@@@@@@@@Oo`***`..,...........,O@OOO@@@@@@@@@@@@....,[ooOOOooOOOOOOoOO^*..*O@OOOOO@@@@@@@@@@@@@@O.=O^..=OOOO\.......      ...     
// ...,O@@@@@@@@^...... ..Oo*=@@@@@O.     .....=@@@@@@@@@@@Oo^*****o...,\`...........[@@@@@@OO@@@@@@\.........*oooOOOOOOoo]****O@OOOOO@@@@@@@@@@@@@@@.*o`..oOOOOO^......      ......  
// ../@@@@@@@@@@^...*.  .=O^*=@@@@@/.     .....=@@@@@@@@@@Oo^*****.=\*..=Oo`...........,O@@@@@@@@OOOOOO`.....,oo[*..=oOOO/`****O@OOOO@@@@@@@@@@@@@@@@^.*...OOOOOOo.......      .......
// ,O@O@@@@@@@@O`.**.   .o/**=@@@@@^      .....=@@@@@@@@@O`****....OO^***OO^******........\@@@@@OOO**=OOO]]oo[*.....//[.*******=@@OO@@@@@@@@@@@@@@@@@O.....OOOOOOO^..*................
// @@OO@@@@@@@@O**/.  ../o***=@@@@O.      .....=O@@@@@@@O^****..*/ooo`**=oO^******..........\@@@OOOOoooOOOOO^.............******@@@@@@@@@@@@@@@@@@@@@@^...,OOOOOOOo..*................
// OOOOO@@@@@@@/*[...]OOO/***=@@@@^      ......=O@@@@@@Oo******/o********\^*****..............,OOO@O`......,OOOO`...........****O@@@@@@@@@@@@@@@@@@@@@O`..=OOOOOOOO^..*...............
